* SPICE NETLIST
***************************************

.SUBCKT Cnt_Active_Auto_10_1
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Cnt_Active_Auto_2_1
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Half_Adder Vdd Gnd Sum Carry A B
** N=13 EP=6 IP=8 FDC=17
M0 3 B Gnd Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=3.375e-13 AS=5.25e-13 PD=1.65e-06 PS=2.9e-06 $X=-4782 $Y=4257 $D=1
M1 Gnd A 3 Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=2.8125e-13 AS=3.375e-13 PD=1.5e-06 PS=1.65e-06 $X=-3632 $Y=4257 $D=1
M2 4 A Gnd Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=1.875e-13 AS=2.8125e-13 PD=1.25e-06 PS=1.5e-06 $X=-2632 $Y=4257 $D=1
M3 Sum B 4 Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=5.0625e-13 AS=1.875e-13 PD=2.1e-06 PS=1.25e-06 $X=-1882 $Y=4257 $D=1
M4 Gnd 3 Sum Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=5.25e-13 AS=5.0625e-13 PD=2.9e-06 PS=2.1e-06 $X=-282 $Y=4257 $D=1
M5 6 A Gnd Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=3.375e-13 AS=5.625e-13 PD=1.65e-06 PS=3e-06 $X=10923 $Y=4291 $D=1
M6 7 B 6 Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=4.875e-13 AS=3.375e-13 PD=2.8e-06 PS=1.65e-06 $X=12073 $Y=4291 $D=1
M7 Gnd 7 Carry Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=5.625e-13 AS=5.625e-13 PD=3e-06 PS=3e-06 $X=20288 $Y=4291 $D=1
M8 9 B 3 Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=5.625e-13 AS=9.375e-13 PD=2.15e-06 PS=4e-06 $X=-4782 $Y=8507 $D=2
M9 Vdd A 9 Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=5.3125e-13 AS=5.625e-13 PD=2.1e-06 PS=2.15e-06 $X=-3632 $Y=8507 $D=2
M10 10 A Vdd Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=3.125e-13 AS=5.3125e-13 PD=1.75e-06 PS=2.1e-06 $X=-2532 $Y=8507 $D=2
M11 Sum 3 10 Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=5.59375e-13 AS=3.125e-13 PD=2.145e-06 PS=1.75e-06 $X=-1782 $Y=8507 $D=2
M12 11 3 Sum Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=3.15625e-13 AS=5.59375e-13 PD=1.755e-06 PS=2.145e-06 $X=-637 $Y=8507 $D=2
M13 Vdd B 11 Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=8.125e-13 AS=3.15625e-13 PD=3.8e-06 PS=1.755e-06 $X=118 $Y=8507 $D=2
M14 7 A Vdd Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=4.6875e-13 AS=9.375e-13 PD=2e-06 PS=4e-06 $X=10923 $Y=8541 $D=2
M15 Vdd B 7 Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=8.75e-13 AS=4.6875e-13 PD=3.9e-06 PS=2e-06 $X=11923 $Y=8541 $D=2
M16 Vdd 7 Carry Vdd PMOS25 L=2.5e-07 W=1.25e-06 AD=9.375e-13 AS=9.375e-13 PD=4e-06 PS=4e-06 $X=20288 $Y=8541 $D=2
.ENDS
***************************************
